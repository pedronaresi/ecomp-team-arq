library verilog;
use verilog.vl_types.all;
entity IO_vlg_vec_tst is
end IO_vlg_vec_tst;
