library verilog;
use verilog.vl_types.all;
entity ExtSinal_vlg_vec_tst is
end ExtSinal_vlg_vec_tst;
