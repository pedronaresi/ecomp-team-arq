library verilog;
use verilog.vl_types.all;
entity MemDados_vlg_vec_tst is
end MemDados_vlg_vec_tst;
