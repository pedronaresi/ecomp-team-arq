library verilog;
use verilog.vl_types.all;
entity BancoReg_vlg_vec_tst is
end BancoReg_vlg_vec_tst;
