module DiscoRigido(clock, trilha, setor, saida, reset, clock_hd, clock_auto, OpHD, pronto, dadosLidos);
	input [31:0] trilha, setor, dadosLidos;
	input clock, clock_hd, clock_auto;
	input reset;
	input [1:0]	OpHD; //0 - nada, 1 - realizar leitura, 2 - realizar gravação
	output reg pronto;
	output reg [31:0] saida;
	parameter size = 2**14;
	
	reg [6:0] aux = 0;
	
	reg [31:0] hd [size-1: 0]; //HD[trilha][setor]
	
	initial
	begin: INIT
	
			//SO
			hd[0] = 0; 		//nome
			hd[1] = 1; 		//trilha
			hd[2] = 3000; 	//tamanho
			hd[3] = 1; 		//ativo
			hd[4] = 0; 		//
			
			//Prog 01
			hd[5] = 5; 		//nome
			hd[6] = 2; 		//trilha
			hd[7] = 500; 	//tamanho
			hd[8] = 1; 		//ativo
			hd[9] = 0; 	//
			
			//Prog 02	
			hd[10] = 6;	 	//nome
			hd[11] = 3; 	//trilha
			hd[12] = 500; 	//tamanho
			hd[13] = 1; 	//ativo
			hd[14] = 0; 	//
			
			//Prog 03	
			hd[15] = 7;	 	//nome
			hd[16] = 4; 	//trilha
			hd[17] = 500; 	//tamanho
			hd[18] = 1; 	//ativo
			hd[19] = 0; 	//
			
			//Prog 04	
			hd[20] = 8;	 	//nome
			hd[21] = 5; 	//trilha
			hd[22] = 500; 	//tamanho
			hd[23] = 1; 	//ativo
			hd[24] = 0; 	//
			
			//Prog 05	
			hd[25] = 2;	 	//nome
			hd[26] = 6; 	//trilha
			hd[27] = 500; 	//tamanho
			hd[28] = 1; 	//ativo
			hd[29] = 0; 	//
			
			//Prog 06	
			hd[30] = 3;	 	//nome
			hd[31] = 7; 	//trilha
			hd[32] = 500; 	//tamanho
			hd[33] = 0; 	//ativo
			hd[34] = 0; 	//
			
			//Prog 07	
			hd[35] = 20;	 	//nome
			hd[36] = 8; 	//trilha
			hd[37] = 500; 	//tamanho
			hd[38] = 0; 	//ativo
			hd[39] = 0; 	//
			
			//Prog 08	
			hd[40] = 9;	 	//nome
			hd[41] = 9; 	//trilha
			hd[42] = 500; 	//tamanho
			hd[43] = 0; 	//ativo
			hd[44] = 0; 	//
			
			//Prog 09	
			hd[45] = 14;	 	//nome
			hd[46] = 10; 	//trilha
			hd[47] = 500; 	//tamanho
			hd[48] = 0; 	//ativo
			hd[49] = 0; 	//
			
			//Prog 10	
			hd[50] = 13;	 	//nome
			hd[51] = 11; 	//trilha
			hd[52] = 500; 	//tamanho
			hd[53] = 0; 	//ativo
			hd[54] = 0; 	//
			
			//Prog 11	
			hd[55] = 24;	 	//nome
			hd[56] = 12; 	//trilha
			hd[57] = 500; 	//tamanho
			hd[58] = 0; 	//ativo
			hd[59] = 0; 	//
			
			//Prog 12	
			hd[60] = 21;	 	//nome
			hd[61] = 13; 	//trilha
			hd[62] = 500; 	//tamanho
			hd[63] = 0; 	//ativo
			hd[64] = 0; 	//
			
			//SO

			hd[100] = 32'b011011_00000_10101_0000001010111100;		//LOADI	21,700
			hd[101] = 32'b000101_11000_10101_01111_00000000000;		//MULT	15,24,21
			hd[102] = 32'b011011_00000_11010_0000000011000111;		//LOADI	26,199
			hd[103] = 32'b000001_01111_11010_11010_00000000000;		//ADD	26,15,26
			hd[104] = 32'b011011_00000_11100_0000000011011111;		//LOADI	28,223
			hd[105] = 32'b000001_01111_11100_11100_00000000000;		//ADD	28,15,28
			hd[106] = 32'b011011_00000_11011_0000000011011100;		//LOADI	27,220
			hd[107] = 32'b000001_01111_11011_11011_00000000000;		//ADD	27,15,27
			hd[108] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[109] = 32'b011011_00000_11110_0000010001111100;		//LOADIR	30,_Fim
			hd[110] = 32'b010100_00000000000000001111111001;		//J	main
			hd[111] = 32'b00000000000000000000000000000000;		//LABEL	findProg
			hd[112] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[113] = 32'b011010_11100_10101_0000000000000010;		//STORE	21,2,28
			hd[114] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[115] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[116] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[117] = 32'b011011_00000_10101_0000000000010000;		//LOADI	21,16
			hd[118] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[119] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[120] = 32'b010110_10110_10101_10101_00000000000;		//SLT	21,22,21
			hd[121] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[122] = 32'b010000_10101_00000_0000000001000010;		//BEQ	21,0,_Fim_While0
			hd[123] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[124] = 32'b011011_00000_10111_0000000000000101;		//LOADI	23,5
			hd[125] = 32'b000101_10111_10101_10101_00000000000;		//MULT	21,23,21
			hd[126] = 32'b000010_10101_10101_0000000000000011;		//ADDI	21,21,3
			hd[127] = 32'b100010_00000_10101_10101_00000000000;		//LOADFT	21,0,21
			hd[128] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[129] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[130] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[131] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[132] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[133] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[134] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[135] = 32'b010000_10101_00000_0000000000110111;		//BEQ	21,0,_Else0
			hd[136] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[137] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[138] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[139] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[140] = 32'b011011_00000_10111_0000000000000101;		//LOADI	23,5
			hd[141] = 32'b000101_10111_10101_10101_00000000000;		//MULT	21,23,21
			hd[142] = 32'b100010_00000_10101_10101_00000000000;		//LOADFT	21,0,21
			hd[143] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[144] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[145] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[146] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[147] = 32'b010000_10101_00000_0000000000110100;		//BEQ	21,0,_Else1
			hd[148] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[149] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[150] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[151] = 32'b010100_00000000000000000000110101;		//J	_Fim_If1
			hd[152] = 32'b00000000000000000000000000000000;		//LABEL	_Else1
			hd[153] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If1
			hd[154] = 32'b010100_00000000000000000000111000;		//J	_Fim_If0
			hd[155] = 32'b00000000000000000000000000000000;		//LABEL	_Else0
			hd[156] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If0
			hd[157] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[158] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[159] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[160] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[161] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[162] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[163] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[164] = 32'b011010_11100_10101_0000000000000010;		//STORE	21,2,28
			hd[165] = 32'b010100_00000000000000000000001110;		//J	14
			hd[166] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_While0
			hd[167] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[168] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[169] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[170] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[171] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[172] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[173] = 32'b000011_10110_10101_10101_00000000000;		//SUB	21,22,21
			hd[174] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[175] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[176] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[177] = 32'b00000000000000000000000000000000;		//LABEL	saveRegs
			hd[178] = 32'b011101_01111_10101_0000000000000000;		//MOVE	21,15
			hd[179] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[180] = 32'b011101_11000_10101_0000000000000000;		//MOVE	21,24
			hd[181] = 32'b011010_11100_10101_0000000000000010;		//STORE	21,2,28
			hd[182] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[183] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[184] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[185] = 32'b011011_00000_10101_0000000011001000;		//LOADI	21,200
			hd[186] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[187] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[188] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[189] = 32'b011010_11100_10101_0000000000000011;		//STORE	21,3,28
			hd[190] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[191] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[192] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[193] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[194] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[195] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[196] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[197] = 32'b011010_10101_00000_0000000000000000;		//STORE	0,0,21
			hd[198] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[199] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[200] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[201] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[202] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[203] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[204] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[205] = 32'b011010_10101_00001_0000000000000000;		//STORE	1,0,21
			hd[206] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[207] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[208] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[209] = 32'b011011_00000_10101_0000000000000010;		//LOADI	21,2
			hd[210] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[211] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[212] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[213] = 32'b011010_10101_00010_0000000000000000;		//STORE	2,0,21
			hd[214] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[215] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[216] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[217] = 32'b011011_00000_10101_0000000000000011;		//LOADI	21,3
			hd[218] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[219] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[220] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[221] = 32'b011010_10101_00011_0000000000000000;		//STORE	3,0,21
			hd[222] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[223] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[224] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[225] = 32'b011011_00000_10101_0000000000000100;		//LOADI	21,4
			hd[226] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[227] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[228] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[229] = 32'b011010_10101_00100_0000000000000000;		//STORE	4,0,21
			hd[230] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[231] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[232] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[233] = 32'b011011_00000_10101_0000000000000101;		//LOADI	21,5
			hd[234] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[235] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[236] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[237] = 32'b011010_10101_00101_0000000000000000;		//STORE	5,0,21
			hd[238] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[239] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[240] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[241] = 32'b011011_00000_10101_0000000000000110;		//LOADI	21,6
			hd[242] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[243] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[244] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[245] = 32'b011010_10101_00110_0000000000000000;		//STORE	6,0,21
			hd[246] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[247] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[248] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[249] = 32'b011011_00000_10101_0000000000000111;		//LOADI	21,7
			hd[250] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[251] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[252] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[253] = 32'b011010_10101_00111_0000000000000000;		//STORE	7,0,21
			hd[254] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[255] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[256] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[257] = 32'b011011_00000_10101_0000000000001000;		//LOADI	21,8
			hd[258] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[259] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[260] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[261] = 32'b011010_10101_01000_0000000000000000;		//STORE	8,0,21
			hd[262] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[263] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[264] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[265] = 32'b011011_00000_10101_0000000000001001;		//LOADI	21,9
			hd[266] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[267] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[268] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[269] = 32'b011010_10101_01001_0000000000000000;		//STORE	9,0,21
			hd[270] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[271] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[272] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[273] = 32'b011011_00000_10101_0000000000001010;		//LOADI	21,10
			hd[274] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[275] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[276] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[277] = 32'b011010_10101_01010_0000000000000000;		//STORE	10,0,21
			hd[278] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[279] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[280] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[281] = 32'b011011_00000_10101_0000000000001011;		//LOADI	21,11
			hd[282] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[283] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[284] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[285] = 32'b011010_10101_01011_0000000000000000;		//STORE	11,0,21
			hd[286] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[287] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[288] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[289] = 32'b011011_00000_10101_0000000000001100;		//LOADI	21,12
			hd[290] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[291] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[292] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[293] = 32'b011010_10101_01100_0000000000000000;		//STORE	12,0,21
			hd[294] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[295] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[296] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[297] = 32'b011011_00000_10101_0000000000001101;		//LOADI	21,13
			hd[298] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[299] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[300] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[301] = 32'b011010_10101_01101_0000000000000000;		//STORE	13,0,21
			hd[302] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[303] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[304] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[305] = 32'b011011_00000_10101_0000000000001110;		//LOADI	21,14
			hd[306] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[307] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[308] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[309] = 32'b011010_10101_01110_0000000000000000;		//STORE	14,0,21
			hd[310] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[311] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[312] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[313] = 32'b011011_00000_10101_0000000000001111;		//LOADI	21,15
			hd[314] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[315] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[316] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[317] = 32'b011010_10101_01111_0000000000000000;		//STORE	15,0,21
			hd[318] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[319] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[320] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[321] = 32'b011011_00000_10101_0000000000010000;		//LOADI	21,16
			hd[322] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[323] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[324] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[325] = 32'b011010_10101_10000_0000000000000000;		//STORE	16,0,21
			hd[326] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[327] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[328] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[329] = 32'b011011_00000_10101_0000000000010001;		//LOADI	21,17
			hd[330] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[331] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[332] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[333] = 32'b011010_10101_10001_0000000000000000;		//STORE	17,0,21
			hd[334] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[335] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[336] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[337] = 32'b011011_00000_10101_0000000000010010;		//LOADI	21,18
			hd[338] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[339] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[340] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[341] = 32'b011010_10101_10010_0000000000000000;		//STORE	18,0,21
			hd[342] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[343] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[344] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[345] = 32'b011011_00000_10101_0000000000010011;		//LOADI	21,19
			hd[346] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[347] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[348] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[349] = 32'b011010_10101_10011_0000000000000000;		//STORE	19,0,21
			hd[350] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[351] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[352] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[353] = 32'b00000000000000000000000000000000;		//LABEL	recoveryRegs
			hd[354] = 32'b011011_00000_10101_0000001010111100;		//LOADI	21,700
			hd[355] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[356] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[357] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[358] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[359] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[360] = 32'b000101_10110_10101_10101_00000000000;		//MULT	21,22,21
			hd[361] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[362] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[363] = 32'b011011_00000_10101_0000000011001000;		//LOADI	21,200
			hd[364] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[365] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[366] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[367] = 32'b011010_11100_10101_0000000000000010;		//STORE	21,2,28
			hd[368] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[369] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[370] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[371] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[372] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[373] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[374] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[375] = 32'b011001_10101_00000_0000000000000000;		//LOAD	0,0,21
			hd[376] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[377] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[378] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[379] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[380] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[381] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[382] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[383] = 32'b011001_10101_00001_0000000000000000;		//LOAD	1,0,21
			hd[384] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[385] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[386] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[387] = 32'b011011_00000_10101_0000000000000010;		//LOADI	21,2
			hd[388] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[389] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[390] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[391] = 32'b011001_10101_00010_0000000000000000;		//LOAD	2,0,21
			hd[392] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[393] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[394] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[395] = 32'b011011_00000_10101_0000000000000011;		//LOADI	21,3
			hd[396] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[397] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[398] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[399] = 32'b011001_10101_00011_0000000000000000;		//LOAD	3,0,21
			hd[400] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[401] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[402] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[403] = 32'b011011_00000_10101_0000000000000100;		//LOADI	21,4
			hd[404] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[405] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[406] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[407] = 32'b011001_10101_00100_0000000000000000;		//LOAD	4,0,21
			hd[408] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[409] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[410] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[411] = 32'b011011_00000_10101_0000000000000101;		//LOADI	21,5
			hd[412] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[413] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[414] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[415] = 32'b011001_10101_00101_0000000000000000;		//LOAD	5,0,21
			hd[416] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[417] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[418] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[419] = 32'b011011_00000_10101_0000000000000110;		//LOADI	21,6
			hd[420] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[421] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[422] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[423] = 32'b011001_10101_00110_0000000000000000;		//LOAD	6,0,21
			hd[424] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[425] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[426] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[427] = 32'b011011_00000_10101_0000000000000111;		//LOADI	21,7
			hd[428] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[429] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[430] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[431] = 32'b011001_10101_00111_0000000000000000;		//LOAD	7,0,21
			hd[432] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[433] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[434] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[435] = 32'b011011_00000_10101_0000000000001000;		//LOADI	21,8
			hd[436] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[437] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[438] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[439] = 32'b011001_10101_01000_0000000000000000;		//LOAD	8,0,21
			hd[440] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[441] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[442] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[443] = 32'b011011_00000_10101_0000000000001001;		//LOADI	21,9
			hd[444] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[445] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[446] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[447] = 32'b011001_10101_01001_0000000000000000;		//LOAD	9,0,21
			hd[448] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[449] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[450] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[451] = 32'b011011_00000_10101_0000000000001010;		//LOADI	21,10
			hd[452] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[453] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[454] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[455] = 32'b011001_10101_01010_0000000000000000;		//LOAD	10,0,21
			hd[456] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[457] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[458] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[459] = 32'b011011_00000_10101_0000000000001011;		//LOADI	21,11
			hd[460] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[461] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[462] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[463] = 32'b011001_10101_01011_0000000000000000;		//LOAD	11,0,21
			hd[464] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[465] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[466] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[467] = 32'b011011_00000_10101_0000000000001100;		//LOADI	21,12
			hd[468] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[469] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[470] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[471] = 32'b011001_10101_01100_0000000000000000;		//LOAD	12,0,21
			hd[472] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[473] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[474] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[475] = 32'b011011_00000_10101_0000000000001101;		//LOADI	21,13
			hd[476] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[477] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[478] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[479] = 32'b011001_10101_01101_0000000000000000;		//LOAD	13,0,21
			hd[480] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[481] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[482] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[483] = 32'b011011_00000_10101_0000000000001110;		//LOADI	21,14
			hd[484] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[485] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[486] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[487] = 32'b011001_10101_01110_0000000000000000;		//LOAD	14,0,21
			hd[488] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[489] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[490] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[491] = 32'b011011_00000_10101_0000000000001111;		//LOADI	21,15
			hd[492] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[493] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[494] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[495] = 32'b011001_10101_01111_0000000000000000;		//LOAD	15,0,21
			hd[496] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[497] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[498] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[499] = 32'b011011_00000_10101_0000000000010000;		//LOADI	21,16
			hd[500] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[501] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[502] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[503] = 32'b011001_10101_10000_0000000000000000;		//LOAD	16,0,21
			hd[504] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[505] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[506] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[507] = 32'b011011_00000_10101_0000000000010001;		//LOADI	21,17
			hd[508] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[509] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[510] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[511] = 32'b011001_10101_10001_0000000000000000;		//LOAD	17,0,21
			hd[512] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[513] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[514] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[515] = 32'b011011_00000_10101_0000000000010010;		//LOADI	21,18
			hd[516] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[517] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[518] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[519] = 32'b011001_10101_10010_0000000000000000;		//LOAD	18,0,21
			hd[520] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[521] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[522] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[523] = 32'b011011_00000_10101_0000000000010011;		//LOADI	21,19
			hd[524] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[525] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[526] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[527] = 32'b011001_10101_10011_0000000000000000;		//LOAD	19,0,21
			hd[528] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[529] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[530] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[531] = 32'b00000000000000000000000000000000;		//LABEL	execProg
			hd[532] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[533] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[534] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[535] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[536] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[537] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[538] = 32'b000011_10110_10101_10101_00000000000;		//SUB	21,22,21
			hd[539] = 32'b011010_11100_10101_0000000000000110;		//STORE	21,6,28
			hd[540] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[541] = 32'b011010_11100_10101_0000000000000101;		//STORE	21,5,28
			hd[542] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[543] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[544] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[545] = 32'b000010_11100_11100_0000000000000111;		//ADDI	28,28,7
			hd[546] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[547] = 32'b000100_11100_11100_0000000000000111;		//SUBI	28,28,7
			hd[548] = 32'b000010_11100_11100_0000000000000111;		//ADDI	28,28,7
			hd[549] = 32'b010101_00000000000000000000001011;		//JAL	findProg
			hd[550] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[551] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[552] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[553] = 32'b000100_11100_11100_0000000000000111;		//SUBI	28,28,7
			hd[554] = 32'b011010_11100_10101_0000000000000011;		//STORE	21,3,28
			hd[555] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[556] = 32'b100000_00000_10101_0000000000000010;		//OUT	2,21
			hd[557] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[558] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[559] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[560] = 32'b011001_11100_10101_0000000000000110;		//LOAD	21,6,28
			hd[561] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[562] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[563] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[564] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[565] = 32'b010000_10101_00000_0000000111011100;		//BEQ	21,0,_Else2
			hd[566] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[567] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[568] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[569] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[570] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[571] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[572] = 32'b000011_10110_10101_10101_00000000000;		//SUB	21,22,21
			hd[573] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[574] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[575] = 32'b010100_00000000000000001000101000;		//J	_Fim_If2
			hd[576] = 32'b00000000000000000000000000000000;		//LABEL	_Else2
			hd[577] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[578] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[579] = 32'b000010_11100_11100_0000000000000111;		//ADDI	28,28,7
			hd[580] = 32'b010101_00000000000000000001001101;		//JAL	saveRegs
			hd[581] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[582] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[583] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[584] = 32'b000100_11100_11100_0000000000000111;		//SUBI	28,28,7
			hd[585] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[586] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[587] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[588] = 32'b000010_11100_11100_0000000000000111;		//ADDI	28,28,7
			hd[589] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[590] = 32'b000100_11100_11100_0000000000000111;		//SUBI	28,28,7
			hd[591] = 32'b000010_11100_11100_0000000000000111;		//ADDI	28,28,7
			hd[592] = 32'b010101_00000000000000000011111101;		//JAL	recoveryRegs
			hd[593] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[594] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[595] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[596] = 32'b000100_11100_11100_0000000000000111;		//SUBI	28,28,7
			hd[597] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[598] = 32'b011101_10101_11000_0000000000000000;		//MOVE	24,21
			hd[599] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[600] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[601] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[602] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[603] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[604] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[605] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[606] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[607] = 32'b010000_10101_00000_0000001000000100;		//BEQ	21,0,_Else3
			hd[608] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[609] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[610] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[611] = 32'b011011_00000_10110_0000000111110100;		//LOADI	22,500
			hd[612] = 32'b000101_10110_10101_10101_00000000000;		//MULT	21,22,21
			hd[613] = 32'b000010_10101_10101_0000100111000100;		//ADDI	21,21,2500
			hd[614] = 32'b100110_10101_11001_0000000000000000;		//JALR	25,21
			hd[615] = 32'b010100_00000000000000001000001001;		//J	_Fim_If3
			hd[616] = 32'b00000000000000000000000000000000;		//LABEL	_Else3
			hd[617] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[618] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[619] = 32'b000010_01010_01010_0000000000000001;		//ADDI	10,10,1
			hd[620] = 32'b100110_01010_11001_0000000000000000;		//JALR	25,10
			hd[621] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If3
			hd[622] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[623] = 32'b011010_11100_10101_0000000000000101;		//STORE	21,5,28
			hd[624] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[625] = 32'b011101_10101_11101_0000000000000000;		//MOVE	29,21
			hd[626] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[627] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[628] = 32'b000010_11100_11100_0000000000000111;		//ADDI	28,28,7
			hd[629] = 32'b010101_00000000000000000001001101;		//JAL	saveRegs
			hd[630] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[631] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[632] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[633] = 32'b000100_11100_11100_0000000000000111;		//SUBI	28,28,7
			hd[634] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[635] = 32'b011101_10101_11000_0000000000000000;		//MOVE	24,21
			hd[636] = 32'b011011_00000_10101_0000001010111100;		//LOADI	21,700
			hd[637] = 32'b000101_11000_10101_01111_00000000000;		//MULT	15,24,21
			hd[638] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[639] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[640] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[641] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[642] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[643] = 32'b000010_11100_11100_0000000000000111;		//ADDI	28,28,7
			hd[644] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[645] = 32'b000100_11100_11100_0000000000000111;		//SUBI	28,28,7
			hd[646] = 32'b000010_11100_11100_0000000000000111;		//ADDI	28,28,7
			hd[647] = 32'b010101_00000000000000000011111101;		//JAL	recoveryRegs
			hd[648] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[649] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[650] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[651] = 32'b000100_11100_11100_0000000000000111;		//SUBI	28,28,7
			hd[652] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If2
			hd[653] = 32'b011001_11100_10101_0000000000000101;		//LOAD	21,5,28
			hd[654] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[655] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[656] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[657] = 32'b00000000000000000000000000000000;		//LABEL	execUmProg
			hd[658] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[659] = 32'b011101_10101_11101_0000000000000000;		//MOVE	29,21
			hd[660] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[661] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[662] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[663] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[664] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[665] = 32'b000010_11100_11100_0000000000000010;		//ADDI	28,28,2
			hd[666] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[667] = 32'b000100_11100_11100_0000000000000010;		//SUBI	28,28,2
			hd[668] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[669] = 32'b000010_11100_11100_0000000000000010;		//ADDI	28,28,2
			hd[670] = 32'b011010_11100_10101_0000000000000010;		//STORE	21,2,28
			hd[671] = 32'b000100_11100_11100_0000000000000010;		//SUBI	28,28,2
			hd[672] = 32'b000010_11100_11100_0000000000000010;		//ADDI	28,28,2
			hd[673] = 32'b010101_00000000000000000110101111;		//JAL	execProg
			hd[674] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[675] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[676] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[677] = 32'b000100_11100_11100_0000000000000010;		//SUBI	28,28,2
			hd[678] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[679] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[680] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[681] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[682] = 32'b00000000000000000000000000000000;		//LABEL	execNProg
			hd[683] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[684] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[685] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[686] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[687] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[688] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[689] = 32'b000011_10110_10101_10101_00000000000;		//SUB	21,22,21
			hd[690] = 32'b011010_11100_10101_0000000000100010;		//STORE	21,34,28
			hd[691] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[692] = 32'b011010_11100_10101_0000000000100001;		//STORE	21,33,28
			hd[693] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[694] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[695] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[696] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[697] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[698] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[699] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[700] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[701] = 32'b010110_10110_10101_10101_00000000000;		//SLT	21,22,21
			hd[702] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[703] = 32'b010000_10101_00000_0000001001111101;		//BEQ	21,0,_Fim_While1
			hd[704] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[705] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[706] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[707] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[708] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[709] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[710] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[711] = 32'b011010_10111_10110_0000000000000010;		//STORE	22,2,23
			hd[712] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[713] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[714] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[715] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[716] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[717] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[718] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[719] = 32'b011010_10111_10110_0000000000001100;		//STORE	22,12,23
			hd[720] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[721] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[722] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[723] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[724] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[725] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[726] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[727] = 32'b011010_10111_10110_0000000000010110;		//STORE	22,22,23
			hd[728] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[729] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[730] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[731] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[732] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[733] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[734] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[735] = 32'b011010_11100_10101_0000000000100001;		//STORE	21,33,28
			hd[736] = 32'b010100_00000000000000001001010011;		//J	595
			hd[737] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_While1
			hd[738] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[739] = 32'b011010_11100_10101_0000000000100001;		//STORE	21,33,28
			hd[740] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[741] = 32'b011010_11100_10101_0000000000100000;		//STORE	21,32,28
			hd[742] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[743] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[744] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[745] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[746] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[747] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[748] = 32'b010110_10110_10101_10101_00000000000;		//SLT	21,22,21
			hd[749] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[750] = 32'b010000_10101_00000_0000001010011110;		//BEQ	21,0,_Fim_While2
			hd[751] = 32'b011001_11100_10101_0000000000100000;		//LOAD	21,32,28
			hd[752] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[753] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[754] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[755] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[756] = 32'b011001_10111_10101_0000000000001100;		//LOAD	21,12,23
			hd[757] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[758] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[759] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[760] = 32'b011010_11100_10101_0000000000100000;		//STORE	21,32,28
			hd[761] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[762] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[763] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[764] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[765] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[766] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[767] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[768] = 32'b011010_11100_10101_0000000000100001;		//STORE	21,33,28
			hd[769] = 32'b010100_00000000000000001010000010;		//J	642
			hd[770] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_While2
			hd[771] = 32'b011001_11100_10101_0000000000100000;		//LOAD	21,32,28
			hd[772] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[773] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[774] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[775] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[776] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[777] = 32'b010111_10110_10101_10101_00000000000;		//SGT	21,22,21
			hd[778] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[779] = 32'b010000_10101_00000_0000001100101011;		//BEQ	21,0,_Fim_While3
			hd[780] = 32'b011001_11100_10101_0000000000100010;		//LOAD	21,34,28
			hd[781] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[782] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[783] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[784] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[785] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[786] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[787] = 32'b011010_11100_10101_0000000000100010;		//STORE	21,34,28
			hd[788] = 32'b011001_11100_10101_0000000000100010;		//LOAD	21,34,28
			hd[789] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[790] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[791] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[792] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[793] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[794] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[795] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[796] = 32'b010000_10101_00000_0000001010111100;		//BEQ	21,0,_Else4
			hd[797] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[798] = 32'b011010_11100_10101_0000000000100010;		//STORE	21,34,28
			hd[799] = 32'b010100_00000000000000001010111101;		//J	_Fim_If4
			hd[800] = 32'b00000000000000000000000000000000;		//LABEL	_Else4
			hd[801] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If4
			hd[802] = 32'b011001_11100_10101_0000000000100010;		//LOAD	21,34,28
			hd[803] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[804] = 32'b011001_10111_10101_0000000000001100;		//LOAD	21,12,23
			hd[805] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[806] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[807] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[808] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[809] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[810] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[811] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[812] = 32'b010000_10101_00000_0000001100000111;		//BEQ	21,0,_Else5
			hd[813] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[814] = 32'b011101_10101_11101_0000000000000000;		//MOVE	29,21
			hd[815] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[816] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[817] = 32'b011001_11100_10101_0000000000100010;		//LOAD	21,34,28
			hd[818] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[819] = 32'b011001_10111_10101_0000000000000010;		//LOAD	21,2,23
			hd[820] = 32'b000010_11100_11100_0000000000100011;		//ADDI	28,28,35
			hd[821] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[822] = 32'b000100_11100_11100_0000000000100011;		//SUBI	28,28,35
			hd[823] = 32'b011001_11100_10101_0000000000100010;		//LOAD	21,34,28
			hd[824] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[825] = 32'b011001_10111_10101_0000000000010110;		//LOAD	21,22,23
			hd[826] = 32'b000010_11100_11100_0000000000100011;		//ADDI	28,28,35
			hd[827] = 32'b011010_11100_10101_0000000000000010;		//STORE	21,2,28
			hd[828] = 32'b000100_11100_11100_0000000000100011;		//SUBI	28,28,35
			hd[829] = 32'b000010_11100_11100_0000000000100011;		//ADDI	28,28,35
			hd[830] = 32'b010101_00000000000000000110101111;		//JAL	execProg
			hd[831] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[832] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[833] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[834] = 32'b000100_11100_11100_0000000000100011;		//SUBI	28,28,35
			hd[835] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[836] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[837] = 32'b011001_11100_10101_0000000000100010;		//LOAD	21,34,28
			hd[838] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[839] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[840] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[841] = 32'b011010_10111_10110_0000000000001100;		//STORE	22,12,23
			hd[842] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[843] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[844] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[845] = 32'b011001_11100_10101_0000000000100010;		//LOAD	21,34,28
			hd[846] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[847] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[848] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[849] = 32'b011010_10111_10110_0000000000010110;		//STORE	22,22,23
			hd[850] = 32'b011001_11100_10101_0000000000100010;		//LOAD	21,34,28
			hd[851] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[852] = 32'b011001_10111_10101_0000000000001100;		//LOAD	21,12,23
			hd[853] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[854] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[855] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[856] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[857] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[858] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[859] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[860] = 32'b010000_10101_00000_0000001100000100;		//BEQ	21,0,_Else6
			hd[861] = 32'b011011_00000_10101_0000000001100100;		//LOADI	21,100
			hd[862] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[863] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[864] = 32'b011001_11100_10101_0000000000100010;		//LOAD	21,34,28
			hd[865] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[866] = 32'b011001_10111_10101_0000000000000010;		//LOAD	21,2,23
			hd[867] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[868] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[869] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[870] = 32'b100000_00000_10101_0000000000000010;		//OUT	2,21
			hd[871] = 32'b010100_00000000000000001100000101;		//J	_Fim_If6
			hd[872] = 32'b00000000000000000000000000000000;		//LABEL	_Else6
			hd[873] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If6
			hd[874] = 32'b010100_00000000000000001100001000;		//J	_Fim_If5
			hd[875] = 32'b00000000000000000000000000000000;		//LABEL	_Else5
			hd[876] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If5
			hd[877] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[878] = 32'b011010_11100_10101_0000000000100001;		//STORE	21,33,28
			hd[879] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[880] = 32'b011010_11100_10101_0000000000100000;		//STORE	21,32,28
			hd[881] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[882] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[883] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[884] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[885] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[886] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[887] = 32'b010110_10110_10101_10101_00000000000;		//SLT	21,22,21
			hd[888] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[889] = 32'b010000_10101_00000_0000001100101001;		//BEQ	21,0,_Fim_While4
			hd[890] = 32'b011001_11100_10101_0000000000100000;		//LOAD	21,32,28
			hd[891] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[892] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[893] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[894] = 32'b000001_10101_11100_10111_00000000000;		//ADD	23,21,28
			hd[895] = 32'b011001_10111_10101_0000000000001100;		//LOAD	21,12,23
			hd[896] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[897] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[898] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[899] = 32'b011010_11100_10101_0000000000100000;		//STORE	21,32,28
			hd[900] = 32'b011001_11100_10101_0000000000100001;		//LOAD	21,33,28
			hd[901] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[902] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[903] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[904] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[905] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[906] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[907] = 32'b011010_11100_10101_0000000000100001;		//STORE	21,33,28
			hd[908] = 32'b010100_00000000000000001100001101;		//J	781
			hd[909] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_While4
			hd[910] = 32'b010100_00000000000000001010011111;		//J	671
			hd[911] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_While3
			hd[912] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[913] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[914] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[915] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[916] = 32'b00000000000000000000000000000000;		//LABEL	renameProg
			hd[917] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[918] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[919] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[920] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[921] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[922] = 32'b000010_11100_11100_0000000000000100;		//ADDI	28,28,4
			hd[923] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[924] = 32'b000100_11100_11100_0000000000000100;		//SUBI	28,28,4
			hd[925] = 32'b000010_11100_11100_0000000000000100;		//ADDI	28,28,4
			hd[926] = 32'b010101_00000000000000000000001011;		//JAL	findProg
			hd[927] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[928] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[929] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[930] = 32'b000100_11100_11100_0000000000000100;		//SUBI	28,28,4
			hd[931] = 32'b011010_11100_10101_0000000000000011;		//STORE	21,3,28
			hd[932] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[933] = 32'b100000_00000_10101_0000000000000010;		//OUT	2,21
			hd[934] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[935] = 32'b011010_11100_10101_0000000000000010;		//STORE	21,2,28
			hd[936] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[937] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[938] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[939] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[940] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[941] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[942] = 32'b011011_00000_10111_0000000000000101;		//LOADI	23,5
			hd[943] = 32'b000101_10111_10110_10110_00000000000;		//MULT	22,23,22
			hd[944] = 32'b100100_10110_00000_10101_00000000000;		//STOREHD	21,0,22
			hd[945] = 32'b100001_10110_00000_10110_00000000000;		//CPHFT	22,0,22
			hd[946] = 32'b011011_00000_10101_0010011100001111;		//LOADI	21,9999
			hd[947] = 32'b100000_00000_10101_0000000000000010;		//OUT	2,21
			hd[948] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[949] = 32'b011011_00000_10111_0000000000000101;		//LOADI	23,5
			hd[950] = 32'b000101_10111_10101_10101_00000000000;		//MULT	21,23,21
			hd[951] = 32'b100010_00000_10101_10101_00000000000;		//LOADFT	21,0,21
			hd[952] = 32'b100000_00000_10101_0000000000000010;		//OUT	2,21
			hd[953] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[954] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[955] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[956] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[957] = 32'b00000000000000000000000000000000;		//LABEL	findEmpty
			hd[958] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[959] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[960] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[961] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[962] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[963] = 32'b011011_00000_10101_0000000000010000;		//LOADI	21,16
			hd[964] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[965] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[966] = 32'b010110_10110_10101_10101_00000000000;		//SLT	21,22,21
			hd[967] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[968] = 32'b010000_10101_00000_0000001110000001;		//BEQ	21,0,_Fim_While5
			hd[969] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[970] = 32'b011011_00000_10111_0000000000000101;		//LOADI	23,5
			hd[971] = 32'b000101_10111_10101_10101_00000000000;		//MULT	21,23,21
			hd[972] = 32'b000010_10101_10101_0000000000000011;		//ADDI	21,21,3
			hd[973] = 32'b100010_00000_10101_10101_00000000000;		//LOADFT	21,0,21
			hd[974] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[975] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[976] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[977] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[978] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[979] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[980] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[981] = 32'b010000_10101_00000_0000001101110110;		//BEQ	21,0,_Else7
			hd[982] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[983] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[984] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[985] = 32'b010100_00000000000000001101110111;		//J	_Fim_If7
			hd[986] = 32'b00000000000000000000000000000000;		//LABEL	_Else7
			hd[987] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If7
			hd[988] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[989] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[990] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[991] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[992] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[993] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[994] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[995] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[996] = 32'b010100_00000000000000001101011100;		//J	860
			hd[997] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_While5
			hd[998] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[999] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1000] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1001] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[1002] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1003] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1004] = 32'b000011_10110_10101_10101_00000000000;		//SUB	21,22,21
			hd[1005] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[1006] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[1007] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[1008] = 32'b00000000000000000000000000000000;		//LABEL	createProg
			hd[1009] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[1010] = 32'b011010_11100_10101_0000000000000100;		//STORE	21,4,28
			hd[1011] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[1012] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1013] = 32'b000010_11100_11100_0000000000000101;		//ADDI	28,28,5
			hd[1014] = 32'b010101_00000000000000001101011001;		//JAL	findEmpty
			hd[1015] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1016] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[1017] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[1018] = 32'b000100_11100_11100_0000000000000101;		//SUBI	28,28,5
			hd[1019] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[1020] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1021] = 32'b100000_00000_10101_0000000000000010;		//OUT	2,21
			hd[1022] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[1023] = 32'b011010_11100_10101_0000000000000010;		//STORE	21,2,28
			hd[1024] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1025] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1026] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1027] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[1028] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1029] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1030] = 32'b011011_00000_10111_0000000000000101;		//LOADI	23,5
			hd[1031] = 32'b000101_10111_10110_10110_00000000000;		//MULT	22,23,22
			hd[1032] = 32'b100100_10110_00000_10101_00000000000;		//STOREHD	21,0,22
			hd[1033] = 32'b100001_10110_00000_10110_00000000000;		//CPHFT	22,0,22
			hd[1034] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[1035] = 32'b011010_11100_10101_0000000000000011;		//STORE	21,3,28
			hd[1036] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1037] = 32'b011011_00000_10111_0000000000000101;		//LOADI	23,5
			hd[1038] = 32'b011011_00000_10110_0000000000000001;		//LOADI	22,1
			hd[1039] = 32'b000101_10111_10101_10101_00000000000;		//MULT	21,23,21
			hd[1040] = 32'b000010_10101_10101_0000000000000011;		//ADDI	21,21,3
			hd[1041] = 32'b100100_10101_00000_10110_00000000000;		//STOREHD	22,0,21
			hd[1042] = 32'b100001_10101_00000_10101_00000000000;		//CPHFT	21,0,21
			hd[1043] = 32'b011001_11100_10101_0000000000000100;		//LOAD	21,4,28
			hd[1044] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1045] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1046] = 32'b011001_11100_10101_0000000000000011;		//LOAD	21,3,28
			hd[1047] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1048] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1049] = 32'b010110_10110_10101_10101_00000000000;		//SLT	21,22,21
			hd[1050] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[1051] = 32'b010000_10101_00000_0000001111011000;		//BEQ	21,0,_Fim_While6
			hd[1052] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[1053] = 32'b011111_00000_10110_0000000000000000;		//IN	22
			hd[1054] = 32'b100111_10110_10101_10111_00000000000;		//ADDU	23,22,21
			hd[1055] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1056] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1057] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1058] = 32'b011001_11100_10101_0000000000000100;		//LOAD	21,4,28
			hd[1059] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1060] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1061] = 32'b000010_10110_10110_0000000000000001;		//ADDI	22,22,1
			hd[1062] = 32'b100100_10101_10110_10111_00000000000;		//STOREHD	23,22,21
			hd[1063] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1064] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1065] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1066] = 32'b011001_11100_10101_0000000000000100;		//LOAD	21,4,28
			hd[1067] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1068] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1069] = 32'b000010_10110_10110_0000000000000001;		//ADDI	22,22,1
			hd[1070] = 32'b011011_00000_10111_0000000111110100;		//LOADI	23,500
			hd[1071] = 32'b000101_10111_10110_10111_00000000000;		//MULT	23,23,22
			hd[1072] = 32'b000010_10111_10111_0000011111010000;		//ADDI	23,23,2000
			hd[1073] = 32'b000001_10111_10101_10111_00000000000;		//ADD	23,23,21
			hd[1074] = 32'b100011_10101_10110_10111_00000000000;		//CPHM	23,22,21
			hd[1075] = 32'b011001_11100_10101_0000000000000100;		//LOAD	21,4,28
			hd[1076] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1077] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1078] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[1079] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1080] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1081] = 32'b000001_10110_10101_10101_00000000000;		//ADD	21,22,21
			hd[1082] = 32'b011010_11100_10101_0000000000000100;		//STORE	21,4,28
			hd[1083] = 32'b010100_00000000000000001110101111;		//J	943
			hd[1084] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_While6
			hd[1085] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[1086] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[1087] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[1088] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[1089] = 32'b00000000000000000000000000000000;		//LABEL	deleteProg
			hd[1090] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[1091] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[1092] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[1093] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1094] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1095] = 32'b000010_11100_11100_0000000000000011;		//ADDI	28,28,3
			hd[1096] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[1097] = 32'b000100_11100_11100_0000000000000011;		//SUBI	28,28,3
			hd[1098] = 32'b000010_11100_11100_0000000000000011;		//ADDI	28,28,3
			hd[1099] = 32'b010101_00000000000000000000001011;		//JAL	findProg
			hd[1100] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1101] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[1102] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[1103] = 32'b000100_11100_11100_0000000000000011;		//SUBI	28,28,3
			hd[1104] = 32'b011010_11100_10101_0000000000000010;		//STORE	21,2,28
			hd[1105] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[1106] = 32'b100000_00000_10101_0000000000000010;		//OUT	2,21
			hd[1107] = 32'b011001_11100_10101_0000000000000010;		//LOAD	21,2,28
			hd[1108] = 32'b011011_00000_10111_0000000000000101;		//LOADI	23,5
			hd[1109] = 32'b000101_10111_10101_10101_00000000000;		//MULT	21,23,21
			hd[1110] = 32'b000010_10101_10101_0000000000000011;		//ADDI	21,21,3
			hd[1111] = 32'b100100_10101_00000_00000_00000000000;		//STOREHD	0,0,21
			hd[1112] = 32'b100001_10101_00000_10101_00000000000;		//CPHFT	21,0,21
			hd[1113] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[1114] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[1115] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[1116] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[1117] = 32'b00000000000000000000000000000000;		//LABEL	main
			hd[1118] = 32'b011011_00000_10101_0000000011001000;		//LOADI	21,200
			hd[1119] = 32'b011010_11011_10101_0000000000000000;		//STORE	21,0,27
			hd[1120] = 32'b011011_00000_10101_0000001010111100;		//LOADI	21,700
			hd[1121] = 32'b011010_11011_10101_0000000000000001;		//STORE	21,1,27
			hd[1122] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[1123] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[1124] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1125] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1126] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1127] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[1128] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1129] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1130] = 32'b010111_10110_10101_10101_00000000000;		//SGT	21,22,21
			hd[1131] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[1132] = 32'b010000_10101_00000_0000010001111000;		//BEQ	21,0,_Fim_While7
			hd[1133] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1134] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1135] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1136] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[1137] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1138] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1139] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[1140] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[1141] = 32'b010000_10101_00000_0000010000011011;		//BEQ	21,0,_Else8
			hd[1142] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[1143] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1144] = 32'b000010_11100_11100_0000000000000010;		//ADDI	28,28,2
			hd[1145] = 32'b010101_00000000000000001000101101;		//JAL	execUmProg
			hd[1146] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1147] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[1148] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[1149] = 32'b000100_11100_11100_0000000000000010;		//SUBI	28,28,2
			hd[1150] = 32'b010100_00000000000000010001110100;		//J	_Fim_If8
			hd[1151] = 32'b00000000000000000000000000000000;		//LABEL	_Else8
			hd[1152] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1153] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1154] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1155] = 32'b011011_00000_10101_0000000000000010;		//LOADI	21,2
			hd[1156] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1157] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1158] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[1159] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[1160] = 32'b010000_10101_00000_0000010000101110;		//BEQ	21,0,_Else9
			hd[1161] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[1162] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1163] = 32'b000010_11100_11100_0000000000000010;		//ADDI	28,28,2
			hd[1164] = 32'b010101_00000000000000001001000110;		//JAL	execNProg
			hd[1165] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1166] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[1167] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[1168] = 32'b000100_11100_11100_0000000000000010;		//SUBI	28,28,2
			hd[1169] = 32'b010100_00000000000000010001110011;		//J	_Fim_If9
			hd[1170] = 32'b00000000000000000000000000000000;		//LABEL	_Else9
			hd[1171] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1172] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1173] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1174] = 32'b011011_00000_10101_0000000000000011;		//LOADI	21,3
			hd[1175] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1176] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1177] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[1178] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[1179] = 32'b010000_10101_00000_0000010001000001;		//BEQ	21,0,_Else10
			hd[1180] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[1181] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1182] = 32'b000010_11100_11100_0000000000000010;		//ADDI	28,28,2
			hd[1183] = 32'b010101_00000000000000001100110000;		//JAL	renameProg
			hd[1184] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1185] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[1186] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[1187] = 32'b000100_11100_11100_0000000000000010;		//SUBI	28,28,2
			hd[1188] = 32'b010100_00000000000000010001110010;		//J	_Fim_If10
			hd[1189] = 32'b00000000000000000000000000000000;		//LABEL	_Else10
			hd[1190] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1191] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1192] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1193] = 32'b011011_00000_10101_0000000000000100;		//LOADI	21,4
			hd[1194] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1195] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1196] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[1197] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[1198] = 32'b010000_10101_00000_0000010001010100;		//BEQ	21,0,_Else11
			hd[1199] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[1200] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1201] = 32'b000010_11100_11100_0000000000000010;		//ADDI	28,28,2
			hd[1202] = 32'b010101_00000000000000001110001100;		//JAL	createProg
			hd[1203] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1204] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[1205] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[1206] = 32'b000100_11100_11100_0000000000000010;		//SUBI	28,28,2
			hd[1207] = 32'b010100_00000000000000010001110001;		//J	_Fim_If11
			hd[1208] = 32'b00000000000000000000000000000000;		//LABEL	_Else11
			hd[1209] = 32'b011001_11100_10101_0000000000000001;		//LOAD	21,1,28
			hd[1210] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1211] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1212] = 32'b011011_00000_10101_0000000000000101;		//LOADI	21,5
			hd[1213] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1214] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1215] = 32'b011000_10110_10101_10101_00000000000;		//SET	21,22,21
			hd[1216] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[1217] = 32'b010000_10101_00000_0000010001100111;		//BEQ	21,0,_Else12
			hd[1218] = 32'b011010_11010_11110_0000000000000000;		//STORE	30,0,26
			hd[1219] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1220] = 32'b000010_11100_11100_0000000000000010;		//ADDI	28,28,2
			hd[1221] = 32'b010101_00000000000000001111011101;		//JAL	deleteProg
			hd[1222] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1223] = 32'b011001_11010_11110_0000000000000000;		//LOAD	30,0,26
			hd[1224] = 32'b011001_11100_10101_0000000000000000;		//LOAD	21,0,28
			hd[1225] = 32'b000100_11100_11100_0000000000000010;		//SUBI	28,28,2
			hd[1226] = 32'b010100_00000000000000010001110000;		//J	_Fim_If12
			hd[1227] = 32'b00000000000000000000000000000000;		//LABEL	_Else12
			hd[1228] = 32'b011011_00000_10101_0000000000000000;		//LOADI	21,0
			hd[1229] = 32'b011010_11010_10101_0000000000000000;		//STORE	21,0,26
			hd[1230] = 32'b000100_11010_11010_0000000000000001;		//SUBI	26,26,1
			hd[1231] = 32'b011011_00000_10101_0000000000000001;		//LOADI	21,1
			hd[1232] = 32'b000010_11010_11010_0000000000000001;		//ADDI	26,26,1
			hd[1233] = 32'b011001_11010_10110_0000000000000000;		//LOAD	22,0,26
			hd[1234] = 32'b000011_10110_10101_10101_00000000000;		//SUB	21,22,21
			hd[1235] = 32'b100000_00000_10101_0000000000000010;		//OUT	2,21
			hd[1236] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If12
			hd[1237] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If11
			hd[1238] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If10
			hd[1239] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If9
			hd[1240] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If8
			hd[1241] = 32'b011111_00000_10101_0000000000000000;		//IN	21
			hd[1242] = 32'b011010_11100_10101_0000000000000001;		//STORE	21,1,28
			hd[1243] = 32'b010100_00000000000000010000000000;		//J	1024
			hd[1244] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_While7
			hd[1245] = 32'b011010_11100_10101_0000000000000000;		//STORE	21,0,28
			hd[1246] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[1247] = 32'b010011_11110_00000_00000_00000000000;		//JR	30
			hd[1248] = 32'b00000000000000000000000000000000;		//LABEL	_Fim
			hd[1249] = 32'b111111_00000000000000000000000000;		//HALT	





	


			//Prog 01
			hd[3000] = 32'b011011_00000_00001_0000001010111100;		//LOADI	1,700
			hd[3001] = 32'b000101_11000_00001_01111_00000000000;		//MULT	15,24,1
			hd[3002] = 32'b011011_00000_01100_0000000011000111;		//LOADI	12,199
			hd[3003] = 32'b000001_01111_01100_01100_00000000000;		//ADD	12,15,12
			hd[3004] = 32'b011011_00000_01110_0000000011011101;		//LOADI	14,221
			hd[3005] = 32'b000001_01111_01110_01110_00000000000;		//ADD	14,15,14
			hd[3006] = 32'b011011_00000_01101_0000000011011100;		//LOADI	13,220
			hd[3007] = 32'b000001_01111_01101_01101_00000000000;		//ADD	13,15,13
			hd[3008] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[3009] = 32'b011011_00000_10000_0000101111101001;		//LOADIR	16,_Fim
			hd[3010] = 32'b010100_00000000000000101111010111;		//J	main
			hd[3011] = 32'b00000000000000000000000000000000;		//LABEL	funcb
			hd[3012] = 32'b011011_00000_00001_0000000000010011;		//LOADI	1,19
			hd[3013] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[3014] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[3015] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[3016] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[3017] = 32'b00000000000000000000000000000000;		//LABEL	func
			hd[3018] = 32'b011011_00000_00001_0000000000010001;		//LOADI	1,17
			hd[3019] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[3020] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[3021] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[3022] = 32'b011010_01100_10000_0000000000000000;		//STORE	16,0,12
			hd[3023] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[3024] = 32'b000010_01110_01110_0000000000000010;		//ADDI	14,14,2
			hd[3025] = 32'b010101_00000000000000101111000011;		//JAL	funcb
			hd[3026] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[3027] = 32'b011001_01100_10000_0000000000000000;		//LOAD	16,0,12
			hd[3028] = 32'b011001_01110_00001_0000000000000000;		//LOAD	1,0,14
			hd[3029] = 32'b000100_01110_01110_0000000000000010;		//SUBI	14,14,2
			hd[3030] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[3031] = 32'b00000000000000000000000000000000;		//LABEL	main
			hd[3032] = 32'b011011_00000_00001_0000000000001111;		//LOADI	1,15
			hd[3033] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[3034] = 32'b011011_00000_00001_0000000000001100;		//LOADI	1,12
			hd[3035] = 32'b011010_01110_00001_0000000000000010;		//STORE	1,2,14
			hd[3036] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[3037] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[3038] = 32'b011010_01100_10000_0000000000000000;		//STORE	16,0,12
			hd[3039] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[3040] = 32'b000010_01110_01110_0000000000000011;		//ADDI	14,14,3
			hd[3041] = 32'b010101_00000000000000101111001001;		//JAL	func
			hd[3042] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[3043] = 32'b011001_01100_10000_0000000000000000;		//LOAD	16,0,12
			hd[3044] = 32'b011001_01110_00001_0000000000000000;		//LOAD	1,0,14
			hd[3045] = 32'b000100_01110_01110_0000000000000011;		//SUBI	14,14,3
			hd[3046] = 32'b011001_01110_00001_0000000000000010;		//LOAD	1,2,14
			hd[3047] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[3048] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[3049] = 32'b00000000000000000000000000000000;		//LABEL	_Fim
			hd[3050] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[3051] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[3052] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[3053] = 32'b111111_00000000000000000000000000;		//HALT	


			
			
			//Prog 02
			hd[3500] = 32'b011011_00000_00001_0000001010111100;		//LOADI	1,700
			hd[3501] = 32'b000101_11000_00001_01111_00000000000;		//MULT	15,24,1
			hd[3502] = 32'b011011_00000_01100_0000000011000111;		//LOADI	12,199
			hd[3503] = 32'b000001_01111_01100_01100_00000000000;		//ADD	12,15,12
			hd[3504] = 32'b011011_00000_01110_0000000011011101;		//LOADI	14,221
			hd[3505] = 32'b000001_01111_01110_01110_00000000000;		//ADD	14,15,14
			hd[3506] = 32'b011011_00000_01101_0000000011011100;		//LOADI	13,220
			hd[3507] = 32'b000001_01111_01101_01101_00000000000;		//ADD	13,15,13
			hd[3508] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[3509] = 32'b011011_00000_10000_0000110111011101;		//LOADIR	16,_Fim
			hd[3510] = 32'b010100_00000000000000110111001011;		//J	main
			hd[3511] = 32'b00000000000000000000000000000000;		//LABEL	funcb
			hd[3512] = 32'b011011_00000_00001_0000000000001001;		//LOADI	1,9
			hd[3513] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[3514] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[3515] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[3516] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[3517] = 32'b00000000000000000000000000000000;		//LABEL	func
			hd[3518] = 32'b011011_00000_00001_0000000000000111;		//LOADI	1,7
			hd[3519] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[3520] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[3521] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[3522] = 32'b011010_01100_10000_0000000000000000;		//STORE	16,0,12
			hd[3523] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[3524] = 32'b000010_01110_01110_0000000000000010;		//ADDI	14,14,2
			hd[3525] = 32'b010101_00000000000000110110110111;		//JAL	funcb
			hd[3526] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[3527] = 32'b011001_01100_10000_0000000000000000;		//LOAD	16,0,12
			hd[3528] = 32'b011001_01110_00001_0000000000000000;		//LOAD	1,0,14
			hd[3529] = 32'b000100_01110_01110_0000000000000010;		//SUBI	14,14,2
			hd[3530] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[3531] = 32'b00000000000000000000000000000000;		//LABEL	main
			hd[3532] = 32'b011011_00000_00001_0000000000000101;		//LOADI	1,5
			hd[3533] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[3534] = 32'b011011_00000_00001_0000000000000010;		//LOADI	1,2
			hd[3535] = 32'b011010_01110_00001_0000000000000010;		//STORE	1,2,14
			hd[3536] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[3537] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[3538] = 32'b011010_01100_10000_0000000000000000;		//STORE	16,0,12
			hd[3539] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[3540] = 32'b000010_01110_01110_0000000000000011;		//ADDI	14,14,3
			hd[3541] = 32'b010101_00000000000000110110111101;		//JAL	func
			hd[3542] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[3543] = 32'b011001_01100_10000_0000000000000000;		//LOAD	16,0,12
			hd[3544] = 32'b011001_01110_00001_0000000000000000;		//LOAD	1,0,14
			hd[3545] = 32'b000100_01110_01110_0000000000000011;		//SUBI	14,14,3
			hd[3546] = 32'b011001_01110_00001_0000000000000010;		//LOAD	1,2,14
			hd[3547] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[3548] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[3549] = 32'b00000000000000000000000000000000;		//LABEL	_Fim
			hd[3550] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[3551] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[3552] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[3553] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[3554] = 32'b111111_00000000000000000000000000;		//HALT	







			//Prog 03
						hd[4000] = 32'b011011_00000_00001_0000001010111100;		//LOADI	1,700
			hd[4001] = 32'b000101_11000_00001_01111_00000000000;		//MULT	15,24,1
			hd[4002] = 32'b011011_00000_01100_0000000011000111;		//LOADI	12,199
			hd[4003] = 32'b000001_01111_01100_01100_00000000000;		//ADD	12,15,12
			hd[4004] = 32'b011011_00000_01110_0000000011011101;		//LOADI	14,221
			hd[4005] = 32'b000001_01111_01110_01110_00000000000;		//ADD	14,15,14
			hd[4006] = 32'b011011_00000_01101_0000000011011100;		//LOADI	13,220
			hd[4007] = 32'b000001_01111_01101_01101_00000000000;		//ADD	13,15,13
			hd[4008] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[4009] = 32'b011011_00000_10000_0000111111010100;		//LOADIR	16,_Fim
			hd[4010] = 32'b010100_00000000000000111111000100;		//J	main
			hd[4011] = 32'b00000000000000000000000000000000;		//LABEL	imprime
			hd[4012] = 32'b011011_00000_00001_0000000000001010;		//LOADI	1,10
			hd[4013] = 32'b011010_01100_00001_0000000000000000;		//STORE	1,0,12
			hd[4014] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[4015] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[4016] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[4017] = 32'b011001_01100_00010_0000000000000000;		//LOAD	2,0,12
			hd[4018] = 32'b010111_00010_00001_00001_00000000000;		//SGT	1,2,1
			hd[4019] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[4020] = 32'b010000_00001_00000_0000111111000000;		//BEQ	1,0,_Fim_While0
			hd[4021] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[4022] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[4023] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[4024] = 32'b011010_01100_00001_0000000000000000;		//STORE	1,0,12
			hd[4025] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[4026] = 32'b011011_00000_00001_0000000000000001;		//LOADI	1,1
			hd[4027] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[4028] = 32'b011001_01100_00010_0000000000000000;		//LOAD	2,0,12
			hd[4029] = 32'b000001_00010_00001_00001_00000000000;		//ADD	1,2,1
			hd[4030] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[4031] = 32'b010100_00000000000000111110101100;		//J	12
			hd[4032] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_While0
			hd[4033] = 32'b011011_00000_00001_0010011100001111;		//LOADI	1,9999
			hd[4034] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[4035] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[4036] = 32'b00000000000000000000000000000000;		//LABEL	main
			hd[4037] = 32'b011111_00000_00001_0000000000000000;		//IN	1
			hd[4038] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[4039] = 32'b011010_01100_10000_0000000000000000;		//STORE	16,0,12
			hd[4040] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[4041] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[4042] = 32'b000010_01110_01110_0000000000000010;		//ADDI	14,14,2
			hd[4043] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[4044] = 32'b000100_01110_01110_0000000000000010;		//SUBI	14,14,2
			hd[4045] = 32'b000010_01110_01110_0000000000000010;		//ADDI	14,14,2
			hd[4046] = 32'b010101_00000000000000111110101011;		//JAL	imprime
			hd[4047] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[4048] = 32'b011001_01100_10000_0000000000000000;		//LOAD	16,0,12
			hd[4049] = 32'b011001_01110_00001_0000000000000000;		//LOAD	1,0,14
			hd[4050] = 32'b000100_01110_01110_0000000000000010;		//SUBI	14,14,2
			hd[4051] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[4052] = 32'b00000000000000000000000000000000;		//LABEL	_Fim
			hd[4053] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[4054] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4055] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[4056] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4057] = 32'b111111_00000000000000000000000000;		//HALT	





		
	
			//Prog 04
			hd[4500] = 32'b011011_00000_00001_0000001010111100;		//LOADI	1,700
			hd[4501] = 32'b000101_11000_00001_01111_00000000000;		//MULT	15,24,1
			hd[4502] = 32'b011011_00000_01100_0000000011000111;		//LOADI	12,199
			hd[4503] = 32'b000001_01111_01100_01100_00000000000;		//ADD	12,15,12
			hd[4504] = 32'b011011_00000_01110_0000000011011101;		//LOADI	14,221
			hd[4505] = 32'b000001_01111_01110_01110_00000000000;		//ADD	14,15,14
			hd[4506] = 32'b011011_00000_01101_0000000011011100;		//LOADI	13,220
			hd[4507] = 32'b000001_01111_01101_01101_00000000000;		//ADD	13,15,13
			hd[4508] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[4509] = 32'b011011_00000_10000_0001000111000111;		//LOADIR	16,_Fim
			hd[4510] = 32'b010100_00000000000001000110101010;		//J	main
			hd[4511] = 32'b00000000000000000000000000000000;		//LABEL	mult
			hd[4512] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[4513] = 32'b011010_01100_00001_0000000000000000;		//STORE	1,0,12
			hd[4514] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[4515] = 32'b011001_01110_00001_0000000000000010;		//LOAD	1,2,14
			hd[4516] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[4517] = 32'b011001_01100_00010_0000000000000000;		//LOAD	2,0,12
			hd[4518] = 32'b000101_00010_00001_00001_00000000000;		//MULT	1,2,1
			hd[4519] = 32'b011010_01110_00001_0000000000000000;		//STORE	1,0,14
			hd[4520] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[4521] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[4522] = 32'b00000000000000000000000000000000;		//LABEL	main
			hd[4523] = 32'b011111_00000_00001_0000000000000000;		//IN	1
			hd[4524] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4525] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4526] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[4527] = 32'b011111_00000_00001_0000000000000000;		//IN	1
			hd[4528] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4529] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4530] = 32'b011010_01110_00001_0000000000000010;		//STORE	1,2,14
			hd[4531] = 32'b011010_01100_10000_0000000000000000;		//STORE	16,0,12
			hd[4532] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[4533] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[4534] = 32'b000010_01110_01110_0000000000000011;		//ADDI	14,14,3
			hd[4535] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[4536] = 32'b000100_01110_01110_0000000000000011;		//SUBI	14,14,3
			hd[4537] = 32'b011001_01110_00001_0000000000000010;		//LOAD	1,2,14
			hd[4538] = 32'b000010_01110_01110_0000000000000011;		//ADDI	14,14,3
			hd[4539] = 32'b011010_01110_00001_0000000000000010;		//STORE	1,2,14
			hd[4540] = 32'b000100_01110_01110_0000000000000011;		//SUBI	14,14,3
			hd[4541] = 32'b000010_01110_01110_0000000000000011;		//ADDI	14,14,3
			hd[4542] = 32'b010101_00000000000001000110011111;		//JAL	mult
			hd[4543] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[4544] = 32'b011001_01100_10000_0000000000000000;		//LOAD	16,0,12
			hd[4545] = 32'b011001_01110_00001_0000000000000000;		//LOAD	1,0,14
			hd[4546] = 32'b000100_01110_01110_0000000000000011;		//SUBI	14,14,3
			hd[4547] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[4548] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4549] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4550] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[4551] = 32'b00000000000000000000000000000000;		//LABEL	_Fim
			hd[4552] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[4553] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4554] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[4555] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[4556] = 32'b111111_00000000000000000000000000;		//HALT	

	




			///Prog 05
			hd[5000] = 32'b011011_00000_00001_0000001010111100;		//LOADI	1,700
			hd[5001] = 32'b000101_11000_00001_01111_00000000000;		//MULT	15,24,1
			hd[5002] = 32'b011011_00000_01100_0000000011000111;		//LOADI	12,199
			hd[5003] = 32'b000001_01111_01100_01100_00000000000;		//ADD	12,15,12
			hd[5004] = 32'b011011_00000_01110_0000000011011101;		//LOADI	14,221
			hd[5005] = 32'b000001_01111_01110_01110_00000000000;		//ADD	14,15,14
			hd[5006] = 32'b011011_00000_01101_0000000011011100;		//LOADI	13,220
			hd[5007] = 32'b000001_01111_01101_01101_00000000000;		//ADD	13,15,13
			hd[5008] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[5009] = 32'b011011_00000_10000_0001001111101001;		//LOADIR	16,_Fim
			hd[5010] = 32'b010100_00000000000001001111000100;		//J	main
			hd[5011] = 32'b00000000000000000000000000000000;		//LABEL	mult
			hd[5012] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[5013] = 32'b011010_01100_00001_0000000000000000;		//STORE	1,0,12
			hd[5014] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[5015] = 32'b011011_00000_00001_0000000000000001;		//LOADI	1,1
			hd[5016] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[5017] = 32'b011001_01100_00010_0000000000000000;		//LOAD	2,0,12
			hd[5018] = 32'b011000_00010_00001_00001_00000000000;		//SET	1,2,1
			hd[5019] = 32'b011011_00000_00000_0000000000000000;		//LOADI	0,0
			hd[5020] = 32'b010000_00001_00000_0001001110100001;		//BEQ	1,0,_Else0
			hd[5021] = 32'b011001_01110_00001_0000000000000010;		//LOAD	1,2,14
			hd[5022] = 32'b011010_01110_00001_0000000000000000;		//STORE	1,0,14
			hd[5023] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[5024] = 32'b010100_00000000000001001110100010;		//J	_Fim_If0
			hd[5025] = 32'b00000000000000000000000000000000;		//LABEL	_Else0
			hd[5026] = 32'b00000000000000000000000000000000;		//LABEL	_Fim_If0
			hd[5027] = 32'b011001_01110_00001_0000000000000010;		//LOAD	1,2,14
			hd[5028] = 32'b011010_01100_00001_0000000000000000;		//STORE	1,0,12
			hd[5029] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[5030] = 32'b011010_01100_10000_0000000000000000;		//STORE	16,0,12
			hd[5031] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[5032] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[5033] = 32'b011010_01100_00001_0000000000000000;		//STORE	1,0,12
			hd[5034] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[5035] = 32'b011011_00000_00001_0000000000000001;		//LOADI	1,1
			hd[5036] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[5037] = 32'b011001_01100_00010_0000000000000000;		//LOAD	2,0,12
			hd[5038] = 32'b000011_00010_00001_00001_00000000000;		//SUB	1,2,1
			hd[5039] = 32'b000010_01110_01110_0000000000000100;		//ADDI	14,14,4
			hd[5040] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[5041] = 32'b000100_01110_01110_0000000000000100;		//SUBI	14,14,4
			hd[5042] = 32'b011001_01110_00001_0000000000000010;		//LOAD	1,2,14
			hd[5043] = 32'b000010_01110_01110_0000000000000100;		//ADDI	14,14,4
			hd[5044] = 32'b011010_01110_00001_0000000000000010;		//STORE	1,2,14
			hd[5045] = 32'b000100_01110_01110_0000000000000100;		//SUBI	14,14,4
			hd[5046] = 32'b000010_01110_01110_0000000000000100;		//ADDI	14,14,4
			hd[5047] = 32'b010101_00000000000001001110010011;		//JAL	mult
			hd[5048] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[5049] = 32'b011001_01100_10000_0000000000000000;		//LOAD	16,0,12
			hd[5050] = 32'b011001_01110_00001_0000000000000000;		//LOAD	1,0,14
			hd[5051] = 32'b000100_01110_01110_0000000000000100;		//SUBI	14,14,4
			hd[5052] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[5053] = 32'b011001_01100_00010_0000000000000000;		//LOAD	2,0,12
			hd[5054] = 32'b000001_00010_00001_00001_00000000000;		//ADD	1,2,1
			hd[5055] = 32'b011010_01110_00001_0000000000000011;		//STORE	1,3,14
			hd[5056] = 32'b011001_01110_00001_0000000000000011;		//LOAD	1,3,14
			hd[5057] = 32'b011010_01110_00001_0000000000000000;		//STORE	1,0,14
			hd[5058] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[5059] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[5060] = 32'b00000000000000000000000000000000;		//LABEL	main
			hd[5061] = 32'b011111_00000_00001_0000000000000000;		//IN	1
			hd[5062] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5063] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5064] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[5065] = 32'b011111_00000_00001_0000000000000000;		//IN	1
			hd[5066] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5067] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5068] = 32'b011010_01110_00001_0000000000000010;		//STORE	1,2,14
			hd[5069] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[5070] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[5071] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5072] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5073] = 32'b011001_01110_00001_0000000000000010;		//LOAD	1,2,14
			hd[5074] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[5075] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5076] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5077] = 32'b011010_01100_10000_0000000000000000;		//STORE	16,0,12
			hd[5078] = 32'b000100_01100_01100_0000000000000001;		//SUBI	12,12,1
			hd[5079] = 32'b011001_01110_00001_0000000000000001;		//LOAD	1,1,14
			hd[5080] = 32'b000010_01110_01110_0000000000000011;		//ADDI	14,14,3
			hd[5081] = 32'b011010_01110_00001_0000000000000001;		//STORE	1,1,14
			hd[5082] = 32'b000100_01110_01110_0000000000000011;		//SUBI	14,14,3
			hd[5083] = 32'b011001_01110_00001_0000000000000010;		//LOAD	1,2,14
			hd[5084] = 32'b000010_01110_01110_0000000000000011;		//ADDI	14,14,3
			hd[5085] = 32'b011010_01110_00001_0000000000000010;		//STORE	1,2,14
			hd[5086] = 32'b000100_01110_01110_0000000000000011;		//SUBI	14,14,3
			hd[5087] = 32'b000010_01110_01110_0000000000000011;		//ADDI	14,14,3
			hd[5088] = 32'b010101_00000000000001001110010011;		//JAL	mult
			hd[5089] = 32'b000010_01100_01100_0000000000000001;		//ADDI	12,12,1
			hd[5090] = 32'b011001_01100_10000_0000000000000000;		//LOAD	16,0,12
			hd[5091] = 32'b011001_01110_00001_0000000000000000;		//LOAD	1,0,14
			hd[5092] = 32'b000100_01110_01110_0000000000000011;		//SUBI	14,14,3
			hd[5093] = 32'b100000_00000_00001_0000000000000010;		//OUT	2,1
			hd[5094] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5095] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5096] = 32'b010011_10000_00000_00000_00000000000;		//JR	16
			hd[5097] = 32'b00000000000000000000000000000000;		//LABEL	_Fim
			hd[5098] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[5099] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5100] = 32'b010011_11001_00000_00000_00000000000;		//JR	25
			hd[5101] = 32'b000000_00000000000000000000000000;		//NOOP	

			hd[5102] = 32'b111111_00000000000000000000000000;		//HALT	





	



	end
	
	
	always @(posedge clock_auto) begin
		
		saida = hd[setor+trilha*(500)*(trilha!=1)+100*(trilha==1)+2000*(trilha>1)];
	end

	
	
	always @(posedge clock) begin
	
		if(OpHD == 2) begin
			hd[setor+trilha*(500)*(trilha!=1)+100*(trilha==1)+2000*(trilha>1)] = dadosLidos;
		end
		
		if(OpHD == 1) begin
			aux = aux + 1;
			if (aux == 2) begin
				pronto = 1;
				aux = 0;
			end
		end
		else if(OpHD == 2) begin
			aux = aux + 1;
			if (aux == 2) begin
				pronto = 1;
				aux = 0;
			end
		end
		else begin 
			pronto = 0;
			aux = 0;
		end 
	end

endmodule	