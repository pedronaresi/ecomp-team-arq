library verilog;
use verilog.vl_types.all;
entity BCD4_vlg_vec_tst is
end BCD4_vlg_vec_tst;
