library verilog;
use verilog.vl_types.all;
entity Processador_vlg_vec_tst is
end Processador_vlg_vec_tst;
