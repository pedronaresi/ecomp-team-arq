library verilog;
use verilog.vl_types.all;
entity Controle_vlg_vec_tst is
end Controle_vlg_vec_tst;
